module risc_cpu (
    input clk, reset    
);
    
endmodule 